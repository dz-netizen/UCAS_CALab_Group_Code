`include "mycpu.h"

//=====================================================================
//  bridge_sram_axi
//  �� CPU �� inst_sram / data_sram ���� ת���� AXI Э��
//  - inst_sram����֧�ֶ�
//  - data_sram��֧�ֶ�/д
//  ���� 4 �� FSM��AR��R��W��B
//=====================================================================

module bridge_sram_axi(
    input  wire          aclk,
    input  wire          aresetn,

    //=================================================================
    // AXI Read Address Channel
    //=================================================================
    output reg  [ 3:0]   arid,        // ������ ID 0=inst,1=data
    output reg  [31:0]   araddr,      // ����ַ
    output reg  [ 7:0]   arlen,       
    output reg  [ 2:0]   arsize,      // �����ݳ��� = log2(8)
    output reg  [ 1:0]   arburst,     // burst type = INCR
    output reg  [ 1:0]   arlock,
    output reg  [ 3:0]   arcache,
    output reg  [ 2:0]   arprot,
    output wire          arvalid,     // �ж�����
    input  wire          arready,     // �������������

    //=================================================================
    // AXI Read Data Channel
    //=================================================================
    input  wire [ 3:0]   rid,         // ���� ID
    input  wire [31:0]   rdata,       // ��������
    input  wire [ 1:0]   rresp,
    input  wire          rlast,       // ���һ�� byte
    input  wire          rvalid,
    output wire          rready,      // ������׼���ý���

    //=================================================================
    // AXI Write Address Channel
    //=================================================================
    output reg  [ 3:0]   awid,        // д��ַ ID = 1
    output reg  [31:0]   awaddr,
    output reg  [ 7:0]   awlen,
    output reg  [ 2:0]   awsize,
    output reg  [ 1:0]   awburst,
    output reg  [ 1:0]   awlock,
    output reg  [ 3:0]   awcache,
    output reg  [ 2:0]   awprot,
    output wire          awvalid,
    input  wire          awready,

    //=================================================================
    // AXI Write Data Channel
    //=================================================================
    output reg  [ 3:0]   wid,         // д ID
    output reg  [31:0]   wdata,
    output reg  [ 3:0]   wstrb,
    output reg           wlast,
    output wire          wvalid,
    input  wire          wready,

    //=================================================================
    // AXI Write Response Channel
    //=================================================================
    input  wire [ 3:0]   bid,
    input  wire [ 1:0]   bresp,
    input  wire          bvalid,
    output wire          bready,

    //=================================================================
    // Inst SRAM interface��������
    //=================================================================
    input  wire          inst_sram_req,
    input  wire          inst_sram_wr,      // ��ԶΪ 0
    input  wire [ 1:0]   inst_sram_size,
    input  wire [31:0]   inst_sram_addr,
    input  wire [ 3:0]   inst_sram_wstrb,
    input  wire [31:0]   inst_sram_wdata,
    output wire          inst_sram_addr_ok, // ��������ַ�ɹ�
    output wire          inst_sram_data_ok, // �յ�������
    output wire [31:0]   inst_sram_rdata,

    //=================================================================
    // Data SRAM interface����/д��
    //=================================================================
    input  wire          data_sram_req,
    input  wire          data_sram_wr,
    input  wire [ 1:0]   data_sram_size,
    input  wire [31:0]   data_sram_addr,
    input  wire [31:0]   data_sram_wdata,
    input  wire [ 3:0]   data_sram_wstrb,
    output wire          data_sram_addr_ok,
    output wire          data_sram_data_ok,
    output wire [31:0]   data_sram_rdata
);

//////////////////////////////////////////////////////////////////////////////////
// �ڲ��źŶ���
//////////////////////////////////////////////////////////////////////////////////

// FSM ״̬������5 bit һ�ȱ���
reg [4:0] ar_current_state, ar_next_state;  // read address
reg [4:0] r_current_state,  r_next_state;   // read data
reg [4:0] w_current_state,  w_next_state;   // write request+data
reg [4:0] b_current_state,  b_next_state;   // write response

// ��Ӧ��������burst ģʽ�¿����ã�
reg [1:0] ar_resp_cnt;
reg [1:0] aw_resp_cnt;
reg [1:0] wd_resp_cnt;

// ������˫���壺buf[0]=inst��buf[1]=data
reg [31:0] buf_rdata [1:0];

// ����д��ͻ
wire read_block;

// ���� rid������ data_ok / inst_ok �ж�
reg [3:0] rid_r;

localparam IDLE = 5'b00001;

//////////////////////////////////////////////////////////////////////////////////
// ������FSM��AR��
//////////////////////////////////////////////////////////////////////////////////

localparam AR_REQ_START = 5'b00010;
localparam AR_REQ_END   = 5'b00100;


// ״̬��ת
always @(posedge aclk) begin
    if (!aresetn)
        ar_current_state <= IDLE;
    else
        ar_current_state <= ar_next_state;
end

// ��һ��״̬
always @(*) begin
    case (ar_current_state)
        IDLE:
            // �������дͬһ����ַ �� ��Ҫ����
            if (read_block)
                ar_next_state = IDLE;

            // inst �� data �Ķ�����
            else if ((data_sram_req & ~data_sram_wr) |
                     (inst_sram_req & ~inst_sram_wr))
                ar_next_state = AR_REQ_START;

            else
                ar_next_state = IDLE;

        AR_REQ_START:
            // ������ handshake �ɹ�
            if (arvalid & arready)
                ar_next_state = AR_REQ_END;
            else
                ar_next_state = AR_REQ_START;

        AR_REQ_END:
            ar_next_state = IDLE;

        default:
            ar_next_state = IDLE;
    endcase
end

assign arvalid = ar_current_state[1];   // ֻ���� START ״̬��������

//////////////////////////////////////////////////////////////////////////////////
// ����Ӧͨ�� FSM��R��
//////////////////////////////////////////////////////////////////////////////////

localparam R_DATA_START = 5'b00010;
localparam R_DATA_END   = 5'b00100;
localparam R_DATA_NEXT   = 5'b01000;
reg con_read_reg;
always @(posedge aclk) begin
    if (!aresetn)
        con_read_reg <=1'b0;
    else if(arvalid & arready & rvalid & rready &rlast&r_current_state[1])
        con_read_reg <= 1'b1;
    else 
        con_read_reg <=1'b0;
end
always @(posedge aclk) begin
    if (!aresetn)
        r_current_state <= IDLE;
    else 
        r_current_state <= r_next_state;
end
reg round;
always @(posedge aclk) begin
    if (!aresetn)
        round <=1'b0;
    else if(r_current_state[1] & arvalid & arready)
        round <=1'b1;
    else if(rvalid & rready)
        round <=1'b0;
end

always @(*) begin
    case (r_current_state)
        IDLE:
            // AR handshake �ɹ���������δ��ɵ� byte
            if (arvalid & arready || |ar_resp_cnt)
                r_next_state = R_DATA_START;
            else
                r_next_state = IDLE;

        R_DATA_START:
            // ���������һ�� beat������������
            if(rvalid & rready & round)
                r_next_state = R_DATA_NEXT;
            else if(arvalid & arready & rvalid & rready &rlast)begin
                r_next_state = R_DATA_START;
            end               
            else if (rvalid & rready & rlast)
                r_next_state = R_DATA_END;
            else
                r_next_state = R_DATA_START;
        R_DATA_NEXT:
             if(rvalid & rready)
                r_next_state = R_DATA_END;
            else
                r_next_state = IDLE;                
        R_DATA_END:
            if(arvalid & arready)
                r_next_state = R_DATA_START;
            else
            r_next_state = IDLE;

        default:begin
            r_next_state = IDLE;
        end
    endcase
end

assign rready = r_current_state[1]|r_current_state[3]; // START ״̬���ն�����

//////////////////////////////////////////////////////////////////////////////////
// д���� + д���� FSM��W��
//////////////////////////////////////////////////////////////////////////////////

localparam W_REQ_START = 5'b00010;  // ��д��ַ��д����
localparam W_ADDR_RESP = 5'b00100;  // �ȴ�д��ַ handshake
localparam W_DATA_RESP = 5'b01000;  // �ȴ�д���� handshake
localparam W_REQ_END   = 5'b10000;  // �ȴ�д��Ӧ B channel

always @(posedge aclk) begin
    if (!aresetn)
        w_current_state <= IDLE;
    else
        w_current_state <= w_next_state;
end

always @(*) begin
    case (w_current_state)
        IDLE:
            if (data_sram_wr)
                w_next_state = W_REQ_START;
            else
                w_next_state = IDLE;

        W_REQ_START:
            // ��ַ������ͬʱ���
            if ((awvalid & awready & wvalid & wready) ||
                ((|aw_resp_cnt)&(|wd_resp_cnt)))
                w_next_state = W_REQ_END;

            // ��ַ�ȳɹ�
            else if (awvalid & awready || |aw_resp_cnt)
                w_next_state = W_ADDR_RESP;

            // �����ȳɹ�
            else if (wvalid & wready || |wd_resp_cnt)
                w_next_state = W_DATA_RESP;

            else
                w_next_state = W_REQ_START;

        W_ADDR_RESP:
            if (wvalid & wready)
                w_next_state = W_REQ_END;
            else
                w_next_state = W_ADDR_RESP;

        W_DATA_RESP:
            if (awvalid & awready)
                w_next_state = W_REQ_END;
            else
                w_next_state = W_DATA_RESP;

        W_REQ_END:
            if (bvalid & bready)
                w_next_state = IDLE;
            else
                w_next_state = W_REQ_END;

        default:
            w_next_state = IDLE;
    endcase
end

assign awvalid = w_current_state[1] | w_current_state[3];
assign wvalid  = w_current_state[1] | w_current_state[2];

//////////////////////////////////////////////////////////////////////////////////
// д��Ӧ FSM��B��
//////////////////////////////////////////////////////////////////////////////////

localparam B_START = 5'b00010;
localparam B_END   = 5'b00100;

always @(posedge aclk) begin
    if (!aresetn)
        b_current_state <= IDLE;
    else
        b_current_state <= b_next_state;
end

always @(*) begin
    case (b_current_state)
        IDLE:
            // �ȴ� W_REQ_END ״̬���� bready
            if (bready)
                b_next_state = B_START;
            else
                b_next_state = IDLE;

        B_START:
            if (bvalid & bready)
                b_next_state = B_END;
            else
                b_next_state = B_START;

        B_END:
            b_next_state = IDLE;

        default:
            b_next_state = IDLE;
    endcase
end

assign bready = w_current_state[4];  // ֻ�� W_REQ_END ״̬����д��Ӧ

//////////////////////////////////////////////////////////////////////////////////
// ����ַ�Ĵ�����ID + ��ַ + size��
//////////////////////////////////////////////////////////////////////////////////

always @(posedge aclk) begin
    if (!aresetn) begin
        arid    <= 0;
        araddr  <= 0;
        arsize  <= 0;
        {arlen, arburst, arlock, arcache, arprot} <= {8'd0,2'b01,1'b0,4'd0,3'd0};
    end
    else if (ar_current_state == IDLE) begin
        // ID ѡ��data ��=1��inst ��=0
        arid   <= {3'b0, data_sram_req & ~data_sram_wr};

        // ��ַѡ��data ����
        araddr <= (data_sram_req & ~data_sram_wr) ? data_sram_addr : inst_sram_addr;

        // size ѡ��
        arsize <= (data_sram_req & ~data_sram_wr) ? 
                  {1'b0, data_sram_size} :
                  {1'b0, inst_sram_size};
    end
end

//////////////////////////////////////////////////////////////////////////////////
// д��ַ�Ĵ���
//////////////////////////////////////////////////////////////////////////////////

always @(posedge aclk) begin
    if (!aresetn) begin
        awaddr <= 0;
        awsize <= 0;
        {awlen, awburst, awlock, awcache, awprot, awid} <=
            {8'd0,2'b01,1'b0,4'd0,3'd0,4'd1};
    end
    else if (w_current_state == IDLE) begin
        awaddr <= data_sram_addr;
        awsize <= {1'b0, data_sram_size};
    end
end

//////////////////////////////////////////////////////////////////////////////////
// д���ݼĴ���
//////////////////////////////////////////////////////////////////////////////////

always @(posedge aclk) begin
    if (!aresetn) begin
        wstrb <= 0;
        wdata <= 0;
        {wid, wlast} <= {4'd1, 1'b1};
    end
    else if (w_current_state == IDLE) begin
        wstrb <= data_sram_wstrb;
        wdata <= data_sram_wdata;
    end
end

//////////////////////////////////////////////////////////////////////////////////
// ��д��ͻ����дͬһ����ַʱ��Ҫ������
//////////////////////////////////////////////////////////////////////////////////

assign read_block =
    (araddr == awaddr) &
    (|w_current_state[4:1]) &
    ~b_current_state[2];

//////////////////////////////////////////////////////////////////////////////////
// �����ݻ��壨���� rid д�룩
//////////////////////////////////////////////////////////////////////////////////

always @(posedge aclk) begin
    if (!aresetn)
        {buf_rdata[1], buf_rdata[0]} <= 64'b0;
    else if (rvalid & rready)
        buf_rdata[rid] <= rdata;
end

assign data_sram_rdata = buf_rdata[1];
assign inst_sram_rdata = buf_rdata[0];

//////////////////////////////////////////////////////////////////////////////////
// addr_ok / data_ok��SRAM �ӿ�����
//////////////////////////////////////////////////////////////////////////////////

assign data_sram_addr_ok =
       arid[0] & arvalid & arready |   // data read ������ַ
       wid[0] & awvalid & awready;     // data write ������ַ

assign data_sram_data_ok =
       rid_r[0] & (r_current_state[2]|con_read_reg)| // data read �յ�����
       bid[0] & bvalid & bready;       // data write �յ���Ӧ

assign inst_sram_addr_ok =
       ~arid[0] & arvalid & arready;   // inst read ������ַ

assign inst_sram_data_ok =
       ~rid_r[0] & (r_current_state[2]|r_current_state[3])| // inst read �յ�����
       ~bid[0] & bvalid & bready;

always @(posedge aclk) begin
    if (!aresetn)
        rid_r <= 0;
    else if (rvalid & rready)
        rid_r <= rid;
end

endmodule
